module sdmoore_tb;
 // Inputs
 logic din;
 logic clk;
 logic reset;

logic [7:0] databits;
 // Outputs
 logic dout;

 // Instantiate the Sequence Detector using Moore FSM
 sdmoore uut (
  .din(din), 
  .clk(clk), 
  .reset(reset), 
  .dout(dout)
 );

// set up the clock
 initial begin
   $dumpfile("dump.vcd");
   $dumpvars(1,uut);
 //  $monitor($time, , ,"clk=%b",clk,,"dout=%b",dout,,"reset=%b",reset,,"din=%b",din);
 clk = 0;
 forever #5 clk = ~clk;
 end 

 initial begin
  // Initialize Inputs
  din = 0; reset =1; databits[7:0] = 8'b01101000;
	#5 reset =0;
	#5;

for (int i = 7 ; i >= 0; i --) begin //Test CORRECT bitstring

	#10 din = databits[i];

end	
	#10;

for (int i = 7; i >= 0; i --) begin //Test CORRECT bitstring

	#10 din = databits[i];

end

	databits[7:0] = 8'b01101001;
	#10;

for (int i = 7; i >= 0; i --) begin //Test WRONG BITSTRING

	#10 din = databits[i];

end

	databits[7:0] = 8'b00110100;
#10;

for (int i = 7; i >= 0; i --) begin //Test WRONG bitstring

	#10 din = databits[i];

end

databits[7:0] = 8'b11010010;


for (int i = 7; i >= 0; i --) begin //Test WRONG Bit string

	#10 din = databits[i];

end
	databits[7:0] = 8'b01101000;
	#10;

for (int i = 7 ; i >= 0; i --) begin //Test CORRECT again

	#10 din = databits[i];

end

	databits[7:0] = 8'b11111111;
	#10;

for (int i = 7; i >= 0; i --) begin //Test WRONG Bit string

	#10 din = databits[i];

end

	databits[7:0] = 8'b10000110;
	#10;

for (int i = 7; i >= 0; i --) begin //Test WRONG Bit string

	#10 din = databits[i];

end



#20 $finish;

end
      

endmodule